module FIR_Filter_L2_Top 
#(
    parameter DATA_IN_WIDTH  = 16,
    parameter DATA_OUT_WIDTH = 64,
    parameter TAP_WIDTH      = 32,
    parameter TAP_COUNT      = 51
)
(
    input wire                               clk,
    input wire                               reset_n,
    input wire   signed [DATA_IN_WIDTH-1:0]  data_in_1,
	 input wire   signed [DATA_IN_WIDTH-1:0]  data_in_2,
    output reg   signed [DATA_OUT_WIDTH-1:0] data_out_1,
	 output reg   signed [DATA_OUT_WIDTH-1:0] data_out_2
);

//input side of diagram
reg [DATA_IN_WIDTH-1:0] data_sum;
assign data_sum = data_in_1 + data_in_2;

// Coefficient values for each tap (to be copied and pasted)
localparam signed [TAP_WIDTH-1:0] H0_taps [0:TAP_COUNT-1] = '{32'b11111111111110000101000100011100, 32'b11111111101101000000010001110011, 32'b11111110110101011110110010000100, 32'b11111101001100100110001111000010, 32'b11111011011001000010101110010000, 32'b11111010111000101110000110111000, 32'b11111100111110010111010100010101, 32'b00000001001011101110100110110101, 32'b00000100111001101000100110000110, 32'b00000101010101100010100111100101, 32'b00000010011000001101001000111111, 32'b11111111001010100000100110100001, 32'b11111111000100011111011111101110, 32'b00000001111101110111111000010001, 32'b00000100001100000000101100011010, 32'b00000010110011110110100011111110, 32'b11111111011011100111010000000100, 32'b11111110011111101100110010101111, 32'b00000001100110100010000111100001, 32'b00000100110011111011100110100011, 32'b00000011001000110110001101011100, 32'b11111101100011000100010101000111, 32'b11111011100011110001010101110010, 32'b00000011010011101001110010101011, 32'b00010001011110111100101000011100, 32'b00011010111110100000001110101110, 32'b00010111100010100111010001011110, 32'b00001010001101001001100110000011, 32'b11111110001010001101000101110100, 32'b11111011100100000011000000011100, 32'b00000000011101000010001100100101, 32'b00000100101110000110100000111010, 32'b00000011100100101110100110111001, 32'b11111111101011011100101000111111, 32'b11111110011011010011001101101110, 32'b00000001000110010010100000101101, 32'b00000011111101111001110010001101, 32'b00000011011011001011111111100001, 32'b00000000010100111100110110111100, 32'b11111110101000000110001000011001, 32'b00000000100010111001101111101100, 32'b00000100001001000010111110000001, 32'b00000101100111111010111100110001, 32'b00000011010011110110001000001100, 32'b11111110111100000101010000001000, 32'b11111011100101000100011110011001, 32'b11111010110111110010101000110100, 32'b11111100001111001011001111010110, 32'b11111110000110010100100000001110, 32'b11111111010111011101110000111000, 32'b11111111111000110010100001001110};

localparam signed [TAP_WIDTH-1:0] H1_taps [0:TAP_COUNT-1] = '{32'b11111111111000110010100001001110, 32'b11111111010111011101110000111000, 32'b11111110000110010100100000001110, 32'b11111100001111001011001111010110, 32'b11111010110111110010101000110100, 32'b11111011100101000100011110011001, 32'b11111110111100000101010000001000, 32'b00000011010011110110001000001100, 32'b00000101100111111010111100110001, 32'b00000100001001000010111110000001, 32'b00000000100010111001101111101100, 32'b11111110101000000110001000011001, 32'b00000000010100111100110110111100, 32'b00000011011011001011111111100001, 32'b00000011111101111001110010001101, 32'b00000001000110010010100000101101, 32'b11111110011011010011001101101110, 32'b11111111101011011100101000111111, 32'b00000011100100101110100110111001, 32'b00000100101110000110100000111010, 32'b00000000011101000010001100100101, 32'b11111011100100000011000000011100, 32'b11111110001010001101000101110100, 32'b00001010001101001001100110000011, 32'b00010111100010100111010001011110, 32'b00011010111110100000001110101110, 32'b00010001011110111100101000011100, 32'b00000011010011101001110010101011, 32'b11111011100011110001010101110010, 32'b11111101100011000100010101000111, 32'b00000011001000110110001101011100, 32'b00000100110011111011100110100011, 32'b00000001100110100010000111100001, 32'b11111110011111101100110010101111, 32'b11111111011011100111010000000100, 32'b00000010110011110110100011111110, 32'b00000100001100000000101100011010, 32'b00000001111101110111111000010001, 32'b11111111000100011111011111101110, 32'b11111111001010100000100110100001, 32'b00000010011000001101001000111111, 32'b00000101010101100010100111100101, 32'b00000100111001101000100110000110, 32'b00000001001011101110100110110101, 32'b11111100111110010111010100010101, 32'b11111010111000101110000110111000, 32'b11111011011001000010101110010000, 32'b11111101001100100110001111000010, 32'b11111110110101011110110010000100, 32'b11111111101101000000010001110011, 32'b11111111111110000101000100011100};

localparam signed [TAP_WIDTH-1:0] H0_H1_taps [0:TAP_COUNT-1] = '{32'b11111111110110110111100101101010, 32'b11111111000100011110000010101011, 32'b11111100111011110011010010010010, 32'b11111001011011110001011110011000, 32'b11110110010000110101010111000100, 32'b11110110011101110010100101010001, 32'b11111011111010011100100100011101, 32'b00000100011111100100101111000001, 32'b00001010100001100011100010110111, 32'b00001001011110100101100101100110, 32'b00000010111011000110111000101011, 32'b11111101110010100110101110111010, 32'b11111111011001011100010110101010, 32'b00000101011001000011110111110010, 32'b00001000001001111010011110100111, 32'b00000011111010001001000100101011, 32'b11111101110110111010011101110010, 32'b11111110001011001001011011101110, 32'b00000101001011010000101110011010, 32'b00001001100010000010000111011101, 32'b00000011100101111000011010000001, 32'b11111001000111000111010101100011, 32'b11111001101101111110011011100110, 32'b00001101100000110011011000101110, 32'b00101001000001100011111001111010, 32'b00110101111101000000011101011100, 32'b00101001000001100011111001111010, 32'b00001101100000110011011000101110, 32'b11111001101101111110011011100110, 32'b11111001000111000111010101100011, 32'b00000011100101111000011010000001, 32'b00001001100010000010000111011101, 32'b00000101001011010000101110011010, 32'b11111110001011001001011011101110, 32'b11111101110110111010011101110010, 32'b00000011111010001001000100101011, 32'b00001000001001111010011110100111, 32'b00000101011001000011110111110010, 32'b11111111011001011100010110101010, 32'b11111101110010100110101110111010, 32'b00000010111011000110111000101011, 32'b00001001011110100101100101100110, 32'b00001010100001100011100010110111, 32'b00000100011111100100101111000001, 32'b11111011111010011100100100011101, 32'b11110110011101110010100101010001, 32'b11110110010000110101010111000100, 32'b11111001011011110001011110011000, 32'b11111100111011110011010010010010, 32'b11111111000100011110000010101011, 32'b11111111110110110111100101101010};


//Data out for sub parallel filters
reg [DATA_OUT_WIDTH-1:0] dataOut_H0;
reg [DATA_OUT_WIDTH-1:0] dataOut_H1;
reg [DATA_OUT_WIDTH-1:0] dataOut_H0H1;

fir_parallel #( .TAPS(H0_taps) ) H0(clk, reset_n, data_in_1, dataOut_H0);
fir_parallel #( .TAPS(H1_taps) ) H1(clk, reset_n, data_in_2, dataOut_H1);
fir_parallel #( .TAPS(H0_H1_taps) ) H0_H1(clk, reset_n, data_sum, dataOut_H0H1);


//output side of diagram:
reg signed [DATA_OUT_WIDTH-1:0] delay;
integer i;
//-----------------------------------------------------------
// Delay Line (for H1)
//-----------------------------------------------------------
always @(posedge clk or negedge reset_n) begin
    if (!reset_n) begin
            delay <= 0;
    end else begin
        // Shift the delay line: new sample enters at delay[0]
        delay <= dataOut_H1;
    end
end


assign data_out_2 = dataOut_H0H1 - dataOut_H1 - dataOut_H0;
assign data_out_1 = dataOut_H0 + delay;

endmodule